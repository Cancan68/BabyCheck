#include "translation.rcp.h"

BITMAPFAMILYEX ID bitmapID_app
BEGIN
  BITMAP "babycheckbw.bmp" BPP 1 COMPRESS DENSITY 1
  BITMAP "babycheck.bmp"   BPP 8 COMPRESS DENSITY 1
  BITMAP "babycheckhr.bmp" BPP 1 COMPRESS DENSITY 2
  BITMAP "babycheckhr.bmp" BPP 8 COMPRESS DENSITY 2
END

ICONFAMILYEX
BEGIN
  BITMAP "babycheckicbw.bmp"  BPP 1 COMPRESS TRANSPARENT 255 255 255
  BITMAP "babycheckic.bmp"    BPP 8 COMPRESS TRANSPARENT 255 255 255 DENSITY 1
  BITMAP "babycheckichr.bmp"  BPP 1 COMPRESS TRANSPARENT 255 255 255 DENSITY 2
  BITMAP "babycheckichr.bmp"  BPP 8 COMPRESS TRANSPARENT 255 255 255 DENSITY 2
END

SMALLICONFAMILYEX
BEGIN
  BITMAP "babychecksmallbw.bmp"   BPP 1 COMPRESS TRANSPARENT 0 255 0
  BITMAP "babychecksmall.bmp"     BPP 8 COMPRESS TRANSPARENT 0 255 0 DENSITY 1
  BITMAP "babychecksmallhr.bmp"   BPP 1 COMPRESS TRANSPARENT 0 255 0 DENSITY 2
  BITMAP "babychecksmallhr.bmp"   BPP 8 COMPRESS TRANSPARENT 0 255 0 DENSITY 2
END

VERSION ID 1 "##VERSION##"
APPLICATIONICONNAME ID 2 "BabyCheck"
APPLICATION ID 3 "CanC"

FORM ID formID_main AT ( 0 0 160 160 )
NOFRAME
MENUID menuID_main
BEGIN
	TITLE "BabyCheck"

        FORMBITMAP 120 105 BITMAP bitmapID_app USABLE
       
        LIST "" ID listID_baby AT (1 20 107 130) USABLE VISIBLEITEMS 10 FONT 0

        BUTTON "MENS" ID buttonID_mes  AT (PREVRIGHT+3 PREVTOP 47 AUTO)
        BUTTON "MOTS" ID buttonID_wor  AT (PREVLEFT PREVBOTTOM+3 47 AUTO)
        BUTTON "ACTION" ID buttonID_action  AT (PREVLEFT PREVBOTTOM+3 47 AUTO)
        BUTTON "SHOTS" ID buttonID_shots  AT (PREVLEFT PREVBOTTOM+3 47 AUTO)
        BUTTON "SYMB" ID buttonID_sym  AT (PREVLEFT PREVBOTTOM+10 47 AUTO)

        BUTTON "NOUV" ID buttonID_new AT (1 140 AUTO AUTO)
        BUTTON "MODI" ID buttonID_ren AT (PREVRIGHT+3 PREVTOP AUTO AUTO)
        BUTTON "SUPP" ID buttonID_sup AT (PREVRIGHT+3 PREVTOP AUTO AUTO)
END

MENU ID menuID_main
BEGIN
        PULLDOWN "BEBE"
        BEGIN
		MENUITEM "NOUVEAU" menuitemID_new "N"
		MENUITEM "MODIFICATION" menuitemID_ren "U"
		MENUITEM "SUPPRIMER" menuitemID_sup "D"
        END
        PULLDOWN "DONNEES"
        BEGIN
                MENUITEM "MENSURATIONS" menuitemID_mes "M"
                MENUITEM "MOTSS" menuitemID_words "W"
                MENUITEM "ACTIONS" menuitemID_action "F"
                MENUITEM "SHOTSS" menuitemID_shots "V"
		MENUITEM SEPARATOR
                MENUITEM "SYMBOLIQUE" menuitemID_symb "S"
        END
        PULLDOWN "INFO"
        BEGIN
                MENUITEM "PREFERENCES" menuitemID_pref "P"
                MENUITEM SEPARATOR
                MENUITEM "INFO" menuitemID_info "I"
                MENUITEM "A_PROPOS" menuitemID_about "A"
        END
END

ALERT ID formID_delete
CONFIRMATION
BEGIN
        TITLE "SUPPRIMER"
        MESSAGE "SUPPRESSION"
        BUTTONS "OK" "CANCEL"
END

FORM ID formID_birth AT(2 4 156 154)
FRAME
MODAL
USABLE
SAVEBEHIND
DEFAULTBTNID buttonID_bircancel
BEGIN
        TITLE "NAISSANCE"

        LABEL "PRENOM"  AUTOID AT (2 20) USABLE FONT 0
        FIELD ID fieldID_firstname AT (PREVRIGHT+3 PREVTOP 100 30) USABLE EDITABLE MULTIPLELINES UNDERLINED AUTOSHIFT MAXCHARS 25 FONT 1

        LABEL "POIDS:"  AUTOID AT (2 PREVBOTTOM+3) USABLE FONT 0
        FIELD ID fieldID_weight AT (PREVRIGHT+3 PREVTOP 30 12) USABLE EDITABLE SINGLELINE MAXCHARS 5 FONT 1
        FIELD ID fieldID_weightu AT (PREVRIGHT+3 PREVTOP 40 12) USABLE NONEDITABLE SINGLELINE MAXCHARS 2 FONT 0

        LABEL "TAILLE:" AUTOID AT (2 PREVBOTTOM+3) USABLE FONT 0
        FIELD ID fieldID_height AT (PREVRIGHT+3 PREVTOP 30 12) USABLE EDITABLE SINGLELINE MAXCHARS 5 FONT 1
        FIELD ID fieldID_heightu AT (PREVRIGHT+3 PREVTOP 30 12) USABLE NONEDITABLE SINGLELINE MAXCHARS 2 FONT 0

	LABEL "DATE_NAI" AUTOID AT (2 PREVBOTTOM+3) USABLE FONT 0
	SELECTORTRIGGER "Mon 00-00-00" ID triggerID_birdate AT(PREVRIGHT+3 PREVTOP AUTO 13) USABLE LEFTANCHOR FONT 1

        LABEL "HEURE" AUTOID AT (2 PREVBOTTOM+3) USABLE FONT 0
	SELECTORTRIGGER "12.00 am" ID triggerID_birtime AT(PREVRIGHT+3 PREVTOP AUTO 13) USABLE LEFTANCHOR FONT 1

        LABEL "SEXE" AUTOID AT (2 PREVBOTTOM+3) USABLE FONT 0
        POPUPTRIGGER "" ID listID_sexet AT (PREVRIGHT+3 PREVTOP 15 13) LEFTANCHOR NOFRAME FONT 0
        POPUPLIST ID listID_sexet listID_sexe
        LIST "M" "F" ID listID_sexe AT (PREVRIGHT+3 PREVTOP 15 13) NONUSABLE DISABLED VISIBLEITEMS 2 FONT 0

        BUTTON "OK" buttonID_birok AT(10 BOTTOM@148 AUTO AUTO) USABLE FONT 0
        BUTTON "CANCEL" buttonID_bircancel AT(PREVRIGHT+4 PREVTOP AUTO AUTO) USABLE FONT 0
END

FORM ID formID_pref AT (30 40 110 81)
FRAME
MODAL
USABLE
SAVEBEHIND
DEFAULTBTNID buttonID_prefcancel
BEGIN
	TITLE "PREFERENCES"

        LABEL "WEIGHTUNIT:" AUTOID AT (2 20) USABLE FONT 0
        POPUPTRIGGER "" ID listID_preftw AT (60 PREVTOP 15 12) LEFTANCHOR NOFRAME FONT 0
	POPUPLIST ID listID_preftw listID_prefw
        LIST "KG" "LB" ID listID_prefw AT (PREVRIGHT+3 PREVTOP 15 12) NONUSABLE DISABLED VISIBLEITEMS 2 FONT 0

        LABEL "HEIGHTUNIT:" AUTOID AT (2 40) USABLE FONT 0
        POPUPTRIGGER "" ID listID_prefth AT (60 PREVTOP 15 12) LEFTANCHOR NOFRAME FONT 0
	POPUPLIST ID listID_prefth listID_prefh
        LIST "CM" "IN" ID listID_prefh AT (PREVRIGHT+3 PREVTOP 15 12) NONUSABLE DISABLED VISIBLEITEMS 2 FONT 0

        BUTTON "OK" buttonID_prefok AT(20 BOTTOM@75 AUTO AUTO) USABLE FONT 0
        BUTTON "CANCEL" buttonID_prefcancel AT(PREVRIGHT+5 PREVTOP AUTO AUTO) USABLE FONT 0
END

FORM ID formID_words AT(0 0 160 160)
FRAME
MODAL
USABLE
SAVEBEHIND
DEFAULTBTNID buttonID_worback
BEGIN
        TITLE "            "

	TABLE ID tableID_words AT (0 15 145 120) ROWS 10 COLUMNS 3 COLUMNWIDTHS 17 40 80

        BUTTON "BACK" buttonID_worback AT(1 PREVBOTTOM+3 AUTO AUTO) USABLE FONT 0
        BUTTON "NOUV" buttonID_wornew AT(PREVRIGHT+3 PREVTOP AUTO AUTO) USABLE FONT 0
        BUTTON "SUPP" buttonID_wordel AT(PREVRIGHT+3 PREVTOP AUTO AUTO) USABLE FONT 0
        BUTTON "Memo" buttonID_wormem AT(PREVRIGHT+3 PREVTOP 32 AUTO) USABLE FONT 0

        SCROLLBAR scrollID_words AT (152 15 7 112) USABLE VALUE 0 MIN 0 MAX 0 PAGESIZE 0
END

FORM ID formID_mesdet AT(2 53 156 105)
FRAME
MODAL
USABLE
SAVEBEHIND
DEFAULTBTNID buttonID_mesdcan
BEGIN
        TITLE "MENSURATIONS"

        LABEL "DATE:" AUTOID AT (20 20) USABLE FONT 0
        SELECTORTRIGGER "Mon 00-00-00" ID triggerID_birdate AT(PREVRIGHT+3 PREVTOP AUTO 13) USABLE LEFTANCHOR FONT 1

        LABEL "POIDS:"  AUTOID AT (20 PREVBOTTOM+3) USABLE FONT 0
        FIELD ID fieldID_weightm AT (PREVRIGHT+3 PREVTOP 30 12) USABLE EDITABLE SINGLELINE MAXCHARS 5 FONT 1
        FIELD ID fieldID_weightu AT (PREVRIGHT+3 PREVTOP 40 12) USABLE NONEDITABLE SINGLELINE MAXCHARS 2 FONT 0

        LABEL "TAILLE:" AUTOID AT (20 PREVBOTTOM+3) USABLE FONT 0
        FIELD ID fieldID_heightm AT (PREVRIGHT+3 PREVTOP 30 12) USABLE EDITABLE SINGLELINE MAXCHARS 5 FONT 1
        FIELD ID fieldID_heightu AT (PREVRIGHT+3 PREVTOP 30 12) USABLE NONEDITABLE SINGLELINE MAXCHARS 2 FONT 0

        LABEL "BMI:" AUTOID AT (20 PREVBOTTOM+3) USABLE FONT 0
        FIELD ID fieldID_bmi AT (PREVRIGHT+3 PREVTOP 30 12) USABLE NONEDITABLE SINGLELINE MAXCHARS 4 FONT 1

        BUTTON "OK" buttonID_mesdok AT(10 PREVBOTTOM+5 AUTO AUTO) USABLE FONT 0
        BUTTON "CANCEL" buttonID_mesdcan AT(PREVRIGHT+4 PREVTOP AUTO AUTO) USABLE FONT 0
        BUTTON "SUPP" buttonID_mesddel AT(PREVRIGHT+4 PREVTOP AUTO AUTO) USABLE FONT 0
END

FORM ID formID_mes AT(0 0 160 160)
FRAME
MODAL
USABLE
SAVEBEHIND
DEFAULTBTNID buttonID_mesback
BEGIN
        TITLE "MENSURATIONS"

        LABEL "DATE"  AUTOID AT (10 13) USABLE FONT 1
        FIELD ID fieldID_weightu AT (55 PREVTOP 40 12) USABLE NONEDITABLE SINGLELINE MAXCHARS 2 FONT 1
        FIELD ID fieldID_heightu AT (88 PREVTOP 30 12) USABLE NONEDITABLE SINGLELINE MAXCHARS 2 FONT 1

        TABLE ID tableID_measur AT (0 PREVBOTTOM+2 110 110) ROWS 10 COLUMNS 3 COLUMNWIDTHS 40 30 30

        SCROLLBAR scrollID_measur AT (111 PREVTOP 7 110) USABLE VALUE 0 MIN 0 MAX 0 PAGESIZE 0

        BUTTON "BACK" buttonID_mesback AT(2 PREVBOTTOM+5 AUTO AUTO) USABLE FONT 0
        BUTTON "NOUV" buttonID_mesnew AT(PREVRIGHT+3 PREVTOP AUTO AUTO) USABLE FONT 0
        BUTTON "Memo" buttonID_mesmem AT(PREVRIGHT+3 PREVTOP AUTO AUTO) USABLE FONT 0

        LABEL "$GRAPH"  AUTOID AT (120 20) USABLE FONT 0
        BUTTON "WEIGHT" buttonID_mesw AT(PREVLEFT PREVBOTTOM+3 38 AUTO) USABLE FONT 0
        BUTTON "HEIGHT" buttonID_mesh AT(PREVLEFT PREVBOTTOM+3 38 AUTO) USABLE FONT 0
        BUTTON "BMI" buttonID_mesbmi AT(PREVLEFT PREVBOTTOM+3 38 AUTO) USABLE FONT 0

END

FORM ID formID_symbol AT(2 53 156 105)
FRAME
MODAL
USABLE
SAVEBEHIND
HELPID stringID_helpsymb
BEGIN
        TITLE "SYMBOLIQUE"

        LABEL "NOMBRE"  AUTOID AT (2 20) USABLE FONT 0
        FIELD ID fieldID_number AT (PREVRIGHT+3 PREVTOP 100 12) USABLE NONEDITABLE SINGLELINE FONT 1

        LABEL "PERIOD"  AUTOID AT (2 35) USABLE FONT 0
        FIELD ID fieldID_period AT (PREVRIGHT+3 PREVTOP 100 12) USABLE NONEDITABLE SINGLELINE FONT 1

        LABEL "SIGNE"  AUTOID AT (2 50) USABLE FONT 0
        FIELD ID fieldID_sign AT (PREVRIGHT+3 PREVTOP 100 12) USABLE NONEDITABLE SINGLELINE FONT 1
        FIELD ID fieldID_signp AT (PREVLEFT PREVBOTTOM+3 100 12) USABLE NONEDITABLE SINGLELINE FONT 1

        BUTTON "OK" buttonID_symok AT(CENTER@78 BOTTOM@103 36 12) USABLE FONT 0
END

FORM ID formID_about AT(2 2 156 156)
FRAME
MODAL
USABLE
SAVEBEHIND
BEGIN
	TITLE "A_PROPOS_T"

        FORMBITMAP 62 15 BITMAP bitmapID_app USABLE

	LABEL "BabyCheck v##VERSION##"	AUTOID AT (CENTER@78 46) USABLE FONT 1
	LABEL "\xA9 Laurent Campredon"	AUTOID AT (CENTER@78 PREVBOTTOM+1) USABLE FONT 0
	LABEL "laurent@campredon.net"		AUTOID AT (CENTER@78 PREVBOTTOM+3) USABLE FONT 1
	LABEL "www.campredon.net"          	AUTOID AT (CENTER@78 PREVBOTTOM+6) USABLE FONT 0
	LABEL "APP_FREEWARE"		AUTOID AT (CENTER@78 PREVBOTTOM+5) USABLE FONT 0

	BUTTON "OK" AUTOID AT(CENTER@78 BOTTOM@150 36 12) USABLE FONT 0
END

FORM ID formID_graph AT(0 0 160 160)
FRAME
MODAL
USABLE
NOSAVEBEHIND
BEGIN
	TITLE "             "

        GADGET ID gadgetID_graph AT (0 15 160 133) USABLE

	BUTTON "OK" buttonID_graphok AT (5 150 AUTO 9) USABLE FONT 0

	PUSHBUTTON "3" ID pushID_3 AT (PREVRIGHT+10 PREVTOP 15 9) USABLE GROUP 1 FONT 0
	PUSHBUTTON "6" ID pushID_6 AT (PREVRIGHT+1 PREVTOP PREVWIDTH 9) USABLE GROUP 1 FONT 0
	PUSHBUTTON "12" ID pushID_12 AT (PREVRIGHT+1 PREVTOP PREVWIDTH 9) USABLE GROUP 1 FONT 0
	PUSHBUTTON "18" ID pushID_18 AT (PREVRIGHT+1 PREVTOP PREVWIDTH 9) USABLE GROUP 1 FONT 0
	PUSHBUTTON "24" ID pushID_24 AT (PREVRIGHT+1 PREVTOP PREVWIDTH 9) USABLE GROUP 1 FONT 0
	PUSHBUTTON "30" ID pushID_30 AT (PREVRIGHT+1 PREVTOP PREVWIDTH 9) USABLE GROUP 1 FONT 0
	PUSHBUTTON "36" ID pushID_36 AT (PREVRIGHT+1 PREVTOP PREVWIDTH 9) USABLE GROUP 1 FONT 0

END

FORM ID formID_shots AT(2 2 156 156)
FRAME
MODAL
USABLE
NOSAVEBEHIND
BEGIN
        TITLE "SHOTSS"

	LABEL "DOCTOR" AUTOID AT (CENTER 13) USABLE FONT 0
        LABEL "DOCTOR2" AUTOID AT (CENTER PREVBOTTOM) USABLE FONT 0

        LABEL "HEB" AUTOID AT (2 44) USABLE FONT 1
        CHECKBOX "" ID checkID_heb1 AT (85 PREVTOP AUTO AUTO) USABLE FONT 0
        CHECKBOX "" ID checkID_heb2 AT (100 PREVTOP AUTO AUTO) USABLE FONT 0
        CHECKBOX "" ID checkID_heb3 AT (115 PREVTOP AUTO AUTO) USABLE FONT 0

        LABEL "DTP" AUTOID AT (2 PREVBOTTOM) USABLE FONT 1
        CHECKBOX "" ID checkID_dtp1 AT (85 PREVTOP AUTO AUTO) USABLE FONT 0
        CHECKBOX "" ID checkID_dtp2 AT (100 PREVTOP AUTO AUTO) USABLE FONT 0
        CHECKBOX "" ID checkID_dtp3 AT (115 PREVTOP AUTO AUTO) USABLE FONT 0
        CHECKBOX "" ID checkID_dtp4 AT (130 PREVTOP AUTO AUTO) USABLE FONT 0

        LABEL "HIB" AUTOID AT (2 PREVBOTTOM) USABLE FONT 1
        CHECKBOX "" ID checkID_hib1 AT (85 PREVTOP AUTO AUTO) USABLE FONT 0
        CHECKBOX "" ID checkID_hib2 AT (100 PREVTOP AUTO AUTO) USABLE FONT 0
        CHECKBOX "" ID checkID_hib3 AT (115 PREVTOP AUTO AUTO) USABLE FONT 0
        CHECKBOX "" ID checkID_hib4 AT (130 PREVTOP AUTO AUTO) USABLE FONT 0

        LABEL "IPV" AUTOID AT (2 PREVBOTTOM) USABLE FONT 1
        CHECKBOX "" ID checkID_ipv1 AT (85 PREVTOP AUTO AUTO) USABLE FONT 0
        CHECKBOX "" ID checkID_ipv2 AT (100 PREVTOP AUTO AUTO) USABLE FONT 0
        CHECKBOX "" ID checkID_ipv3 AT (115 PREVTOP AUTO AUTO) USABLE FONT 0

        LABEL "MMR" AUTOID AT (2 PREVBOTTOM) USABLE FONT 1
        CHECKBOX "" ID checkID_mmr1 AT (85 PREVTOP AUTO AUTO) USABLE FONT 0

        LABEL "VAR" AUTOID AT (2 PREVBOTTOM) USABLE FONT 1
        CHECKBOX "" ID checkID_var1 AT (85 PREVTOP AUTO AUTO) USABLE FONT 0

        LABEL "PCV" AUTOID AT (2 PREVBOTTOM) USABLE FONT 1
        CHECKBOX "" ID checkID_pcv1 AT (85 PREVTOP AUTO AUTO) USABLE FONT 0
        CHECKBOX "" ID checkID_pcv2 AT (100 PREVTOP AUTO AUTO) USABLE FONT 0
        CHECKBOX "" ID checkID_pcv3 AT (115 PREVTOP AUTO AUTO) USABLE FONT 0
        CHECKBOX "" ID checkID_pcv4 AT (130 PREVTOP AUTO AUTO) USABLE FONT 0

        BUTTON "OK" buttonID_shotsok AT (40 PREVBOTTOM+12 AUTO AUTO) USABLE FONT 0
        BUTTON "CANCEL" buttonID_shotscancel AT (PREVRIGHT+3 PREVTOP AUTO AUTO) USABLE FONT 0
END

ALERT ID formID_error
ERROR
BEGIN
        TITLE "ERREUR"
        MESSAGE "^1"
        BUTTONS "OK"
END

ALERT ID formID_info
INFORMATION
BEGIN
        TITLE "INFO"
        MESSAGE "^1"
        BUTTONS "OK"
END

STRING ID stringID_info "AIDE"
STRING ID stringID_selbaby "SELECTBEBE"
STRING ID stringID_birdate "SELECTDATENAISS"
STRING ID stringID_birtime "SELECTTIMENAISS"
STRING ID stringID_wordate "SELECTDATEMOTS"
STRING ID stringID_mesdate "SELECTDATEMESURE"
STRING ID stringID_row "SELECTROW"
STRING ID stringID_romversion "ROMVERSION"
STRING ID stringID_actiondate "SELECTDATEACTION"
STRING ID stringID_shotsdate "SELECTDATESHOTS"
STRING ID stringID_helpsymb "HELPSYMB"
STRING ID stringID_transmemo "TRANSMEMO"
